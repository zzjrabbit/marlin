module main(
    input var clk
);
endmodule
