module veryl_project_Wire (
    input  logic [32-1:0] medium_input ,
    output logic [32-1:0] medium_output
);
    always_comb medium_output = medium_input;
endmodule
//# sourceMappingURL=main.sv.map
