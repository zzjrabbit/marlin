module main(
    input single_input,
    output single_output
);
    assign single_output = single_input;
endmodule
